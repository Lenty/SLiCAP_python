noiseTest
V1 1 0 V value=0 noise = {4*k*T*R_s}
R1 1 3 {R_s}
L1 2 4 {L_s}
C2 3 4 {C_s}
R2 2 0 {R_p}
C1 2 0 {C_p}
R3 3 4 1k
I1 0 2 I value = 0 noise={4*k*T/R_p*(1+f_ell/f)}
.param R_s=1k R_p=1k C_p=1n C_s=1u f_ell=1 L_s=1u
.end
