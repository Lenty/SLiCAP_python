"OptoStage"
.include SLiCAP.lib
C2 1 0 {2*C_pin}
C3 2 0 {C_led}
R3 2 3 {R_led}
R1 4 1 {R_vi}
C1 1 5 {C_f}
R2 5 0 {R_se}
O1 0 1 5 2 AD8610_A0 
F1 0 7 3 6 5m
F2 1 0 6 0 5m
V1 4 0 V value=1 dc=0 dcvar=0 noise=0
.param  C_pin=22p R_vi=51k C_f=4.7p C_led=80p R_led=25 R_se=300 A_0=300k

V2 7 0 V value=0 dc=0 dcvar=0 noise=0
.end
