F.cir
F1 1 2 3 4 myF
R1 1 2 {R_2}
R2 1 3 {R_1}
R3 2 4 {R_1}
R4 1 0 {R_GND}
.model myF F value={A_i*(1+s*tau_z)/(1+s*tau_p)}
.end