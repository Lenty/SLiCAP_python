smallestMatrix
I1 0 1 {I_s}
R1 1 0 {R_s}
.end
