VampBiasTotal
* file: VampBiasTotal.cir
* SLiCAP netlist file
.include SLiCAP.lib
V1 1 0 V dc={V_S} dcvar={(sigma_v*V_S)^2}
R3 1 2 r value={R_a} dcvar={(R_a*sigma_r)^2}
R4 2 0 r value={R_b} dcvar={(R_b*sigma_r)^2}
R6 2 3 r value={R_c} dcvar={(R_c*sigma_r)^2}
R2 out 4 r value={19*R} dcvar={(19*R*sigma_r)^2}
X 4 3 out 0 O_dcvar 
+ sib={I_b*sigma_Ib} 
+ sio={i_off} 
+ svo={v_off} 
+ iib={I_b}
.param R_b={R_a}
.end 
