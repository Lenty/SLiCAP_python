EZ.cir
EZ1 1 2 3 4 myE
R1 1 4 {R_1}
R2 2 3 {R_1}
R3 3 4 {R_2}
R4 1 0 {R_GND}
.model myE EZ value={A_v*(1+s*tau_z)/(1+s*tau_p)} zo={R*(1+s*tau_zz)/(1+s*tau_zp)}
.end