"preamp"
.param R_s=50
R2 2 1 {R_s}
N1 outP 0 1 3
R4 3 outP {R_2}
R3 3 0 {R_3}
E1 outN 0 outP 0 -1
R1 1 outN {R_1}
I1 1 outN {4*k*T/R_1}
I3 3 outP {4*k*T/R_2}
I2 0 3 {4*k*T/R_3}
V1 2 0 {4*k*T*R_s}
.end
