"MOSamp"
.include SLiCAP.lib
V1 1 0 V value = 1
C2 0 out {C_ell}
R1 1 2 {R_s}
R2 0 3 {R_b}
R4 4 out {R_c}
X2 5 0 6 0 CMOS18P W=180n L=180n ID=70n
X5 7 0 8 0 CMOS18P W=180n L=180n ID=35n
X4 5 5 0 0 CMOS18N W=180n L=1u ID=70n
X3 8 0 7 0 CMOS18N W=180n L=180n ID=35n
X8 4 7 0 0 CMOS18N W=3u L=180n ID={I_N}
X7 4 8 0 0 CMOS18P W=5.5u L=180n ID={I_P}
X6 7 5 0 0 CMOS18N W=180n L=1u ID=70n
X1 8 6 2 3 CMOS18ND ID=200n W=180n L=180n
R3 3 4 {R_a}
C1 3 4 {C_c}
.param R_s=1M R_a=9M R_b=1M R_c=1k C_ell=100p C_c={700f} I_P={37n+I_source} I_N={37n+I_sink} I_source=100n I_sink=0
.end
