"Balanced Line Driver"
* Z:\mnt\DATA\SLiCAP\SLiCAP_github\SLiCAP_python\files\examples\balancedAmp\cir\balancedAmp.asc
O1N inN fbN outN 0 OPA627_A0
R2 fbP fbN R value={R_a} noisetemp=0 noiseflow=0 dcvar=0
R3P outP fbP R value={R_b} noisetemp=0 noiseflow=0 dcvar=0
O1P inP fbP outP 0 OPA627_A0
R3N fbN outN R value={R_b} noisetemp=0 noiseflow=0 dcvar=0
C1 outP outN C value={C_d} vinit=0
C2P outP 0 C value={C_c/2} vinit=0
C2N outN 0 C value={C_c/2} vinit=0
V1P scP 0 V value={V_s} dc=0 dcvar=0 noise=0
V1N scN 0 V value=0 dc=0 dcvar=0 noise=0
R1P inP scP R value={R_s} noisetemp=0 noiseflow=0 dcvar=0
R1N inN scN R value={R_s} noisetemp=0 noiseflow=0 dcvar=0
.param R_s=50 R_a=15 R_b=2740 C_d=1n C_c=2n A0=1M
.backanno
.end
