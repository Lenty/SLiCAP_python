"My first RC network"
* Z:\mnt\DATA\SLiCAP\SLiCAP_github\SLiCAP_python\files\examples\myFirstRCnetwork\cir\myFirstRCnetwork.asc
V1 N001 0 V value=1 dc=0 dcvar=0 noise=0
R1 N001 out {R}
C1 out 0 {C}
.param R=1k C={1/(2*pi*R*f_c)} f_c=1k
.backanno
.end
