myFirstVampOPA211bias
XU1 N003 N004 out 0 O_dcvar svo=40u sib=60n sio=30n iib=0
V1 N001 0 V value=0 dc=5 dcvar={(0.0033*5)^2} noise=0
R1 N003 N002 r value=20k dcvar={(0.0033*20k)^2}
R2 out N004 r value=20k dcvar={(0.0033*20k)^2}
R3 N002 N001 r value=1k dcvar={(0.0033*1k)^2}
R4 0 N002 r value=1k dcvar={(0.0033*1k)^2}
.end
