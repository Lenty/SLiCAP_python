defaultParams
Q1 1 1 0 0 QV
.end
