"T circuit -1-"
* Z:\mnt\DATA\SLiCAP\SLiCAP_github\SLiCAP_python\files\examples\balancedCircuits\cir\Tcircuit1.asc
R1 inP C R value={R_a} noisetemp=0 noiseflow=0 dcvar=0
R2 C inN R value={R_b} noisetemp=0 noiseflow=0 dcvar=0
I1 0 inP I value=0 dc=0 dcvar=0 noise=0
I2 0 inN I value=0 dc=0 dcvar=0 noise=0
R3 0 C R value={R_c} noisetemp=0 noiseflow=0 dcvar=0
.backanno
.end
