V.cir
V1 1 2 1
R1 1 3 {R_1}
R2 2 4 {R_1}
R3 3 4 {R_2}
R4 2 0 {R_GND}
.end
