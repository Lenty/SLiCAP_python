"Balanced Line Driver"
* Z:\home\anton\SLiCAP\examples\balancedAmp\cir\balancedAmp.asc
O1N inN fbN outN 0 OPA627_A0
R2 fbP fbN R value=15 noisetemp=0 noiseflow=0 dcvar=0
R3P outP fbP R value=2.74k noisetemp=0 noiseflow=0 dcvar=0
O1P inP fbP outP 0 OPA627_A0
R3N fbN outN R value=2.74k noisetemp=0 noiseflow=0 dcvar=0
C1 outP outN C value=1n vinit=0
C2P outP 0 C value=1n vinit=0
C2N outN 0 C value=1n vinit=0
V1P scP 0 V value=1 dc=0 dcvar=0 noise=0
V1N scN 0 V value=0 dc=0 dcvar=0 noise=0
R1P inP scP R value=50 noisetemp=0 noiseflow=0 dcvar=0
R1N inN scN R value=50 noisetemp=0 noiseflow=0 dcvar=0
.param A0=1M
.backanno
.end
