"Low-pass RL filter"
L1 2 1 {L_a*R}
L2 1 out {L_b*R}
C1 1 0 {C_a/R}
C2 out 0 {C_b/R}
R1 out 0 {R}
.param R=6
V1 2 0 V value=1 dc=0 dcvar=0 noise=0
.end
