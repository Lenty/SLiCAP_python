"AD8610 circuit compensated"
* file: transimpedanceOpampComp.cir
* SLiCAP circuit file
.include SLiCAP.lib
I1 0 1 {I_s}
C1 0 1 {C_s}
R1 1 ell {R_f}
C2 1 ell {C_c}
O1 0 1 ell 0 AD8610
.param 
+ I_s=1 C_s=20p R_f=50k C_c=0
.end
