mosEKVplots
* SLiCAP netlist file
.include SLiCAP.lib
X1 d g s 0 CMOS18P W={W} L={L} ID={I_D}
.param W=220n L=180n
.end
