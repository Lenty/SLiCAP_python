CSresNoise
V1 N001 0 V value=0 dc=0 dcvar=0 noise=0
R1 N001 P001 R value={R_s} noisetemp={T} noiseflow=0 dcvar=0
X1 P001 0 out NM18_noise ID={ID} IG={IG} W={W} L={L}
.param R_s=600 W=54.6u L=180n ID=6.15m IG=0
.end
