"Feedback concept"
* Z:\home\anton\DATA\SLiCAP\Examples\transimpedance\transimpedanceIdeal.asc
C1 N001 0 {C_s}
I1 N001 0 I value={I_s} dc=0 dcvar=0 noise=0
R1 out 0 {R_ell}
C2 out 0 {C_ell}
N1 out 0 N001 0
R2 out N001 {R_f}
.param C_s=20p R_f=100k R_ell=1k C_ell=20p
.backanno
.end
