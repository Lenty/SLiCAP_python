"balanced LPF"
C2 2 1 {C_1}
C3 3 0 {C_2}
.param C_1=2.2n R_1=1.8k
R2 4 2 {R_1}
R3 0 1 {R_1}
R4 2 5 {R_3}
R6 1 3 {R_3}
R5 1 0 {R_2}
C1 5 out {C_2}
N1 out 0 5 3
R1 2 out {R_2}
V1 0 4 1
.end
