"AD8610 circuit"
* file: transimpedanceOpamp.cir
* SLiCAP circuit file
.include SLiCAP.lib
I1 0 1 {I_s}
C1 0 1 {C_s}
R1 1 ell {R_f}
O1 0 1 ell 0 AD8610
.param I_s=1 C_s=20p R_f=50k
.end
