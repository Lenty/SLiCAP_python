Tcircuit1
R1 inP C R value={R_a} noisetemp={T} noiseflow=0 dcvar=0
R2 C inN R value={R_b} noisetemp={T} noiseflow=0 dcvar=0
I2 0 inN I value={I_B} dc=0 dcvar=0 noise={S_B}
I1 0 inP I value={I_A} dc=0 dcvar=0 noise={S_A}
R3 0 C R value={R_c} noisetemp=0 noiseflow=0 dcvar=0
.end
