"LowPassLR"
L1 2 1 {L_a*R}
L2 1 out {L_b*R}
C1 1 0 {C_a/R}
C2 out 0 {C_b/R}
R1 out 0 {R}
V1 2 0 V value={A*s/(s^2+(2*pi*f)^2)} ; cosine, amplitude: A, frequency: f
*V1 2 0 V value={A*2*pi*f/(s^2+(2*pi*f)^2)} ; sine, amplitude: A, frequency: f
.param R=6 C_a=126.6u L_a=150.1u L_b=75.03u C_b=28.13u A=0.5 f=2k
.end
