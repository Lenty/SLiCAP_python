G.cir
G1 1 2 3 4 myG
R1 1 2 {R_2}
R2 1 3 {R_1}
R3 2 4 {R_1}
R4 3 4 {R_3}
R5 1 0 {R_GND}
.model myG G value={A_y*(1+s*tau_z)/(1+s*tau_p)}
.end
